// module header();
//     parameter dwidth_dat = 16;
//     parameter awidth_mem = 12;
//     parameter awidth_reg = 6;
// endmodule


`ifndef _my_incl_vh_
    `define _my_incl_vh_
    // Start of include contents
    `define dwidth_dat 16
    `define awidth_mem 12
    `define awidth_reg 6
    `define inst_start 31
    `define clk_div 125000
    `define dwidth_mat 4
    `define dwidth_dat_user 4
    //`define clk_div 2
`endif
